module mac (
input logic CLK,
input 



);

endmodule 